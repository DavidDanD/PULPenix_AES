`include "../../axi/axi_spi_master/spi_master_fifo.sv"